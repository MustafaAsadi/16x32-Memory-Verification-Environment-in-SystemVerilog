class out_trans;
  logic [31:0] Data_out;
  bit Valid_out;
endclass
